----------------------------------------------
---------------MEMÓRIA ROM--------------------
----------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity rom is
    port 
    (
        clk  : in std_logic;
        addr : in unsigned (7 downto 0);
        data : out unsigned (14 downto 0)
    );
end rom;

architecture a_rom of rom is

    type mem is array (0 to 255) of unsigned (14 downto 0);

    constant conteudo_rom : mem := 
    (
        0	=>	B"0101_00100001_001", 	-- mov r1, #33
        1	=>	B"0101_00000001_010", 	-- mov r2, #1
        2	=>	B"0101_00000001_011", 	-- mov r3, #1
        3	=>	B"0101_00010001_101", 	-- mov r5, #17
        4	=>	B"1000_00000000_000", 	-- mov a, #0
        5	=>	B"0001_00000_010_000", 	-- add a, r2
        6	=>	B"1010_00000_010_000", 	-- mov @r2, a
        7	=>	B"0001_00000_011_000", 	-- add a, r3
        8	=>	B"0110_00000_000_010", 	-- mov r2, a
        9	=>	B"0111_00000000000", 	-- clr c
        10	=>	B"0010_00000_001_000", 	-- subb a, r1
        11	=>	B"1110_000_11111000", 	-- jc inicializa_ram
        12	=>	B"0101_00000010_010", 	-- mov r2, #2
        13	=>	B"1001_00000_010_000", 	-- mov a, @r2
        14	=>	B"0110_00000_000_100", 	-- mov r4, a
        15	=>	B"1000_00000000_000", 	-- mov a, #0
        16	=>	B"0111_00000000000", 	-- clr c
        17	=>	B"0010_00000_100_000", 	-- subb a, r4
        18	=>	B"1110_000_00001000", 	-- jc primo
        19	=>	B"1000_00000000_000", 	-- mov a, #0
        20	=>	B"0001_00000_010_000", 	-- add a, r2
        21	=>	B"0001_00000_011_000", 	-- add a, r3
        22	=>	B"0110_00000_000_010", 	-- mov r2, a
        23	=>	B"0111_00000000000", 	-- clr c
        24	=>	B"0010_00000_101_000", 	-- subb a, r5
        25	=>	B"1110_000_11110011", 	-- jc loop
        26	=>	B"1111_000_00101110", 	-- ajmp fim_loop
        27	=>	B"1000_00000000_000", 	-- mov a, #0
        28	=>	B"0001_00000_100_000", 	-- add a, r4
        29	=>	B"0001_00000_100_000", 	-- add a, r4
        30	=>	B"0110_00000_000_110", 	-- mov r6, a
        31	=>	B"1000_00000000_000", 	-- mov a, #0
        32	=>	B"1010_00000_110_000", 	-- mov @r6, a
        33	=>	B"0001_00000_110_000", 	-- add a, r6
        34	=>	B"0001_00000_100_000", 	-- add a, r4
        35	=>	B"0110_00000_000_110", 	-- mov r6, a
        36	=>	B"0111_00000000000", 	-- clr c
        37	=>	B"0010_00000_001_000", 	-- subb a, r1
        38	=>	B"1110_000_11111000", 	-- jc loop2
        39	=>	B"1000_00000000_000", 	-- mov a, #0
        40	=>	B"0001_00000_010_000", 	-- add a, r2
        41	=>	B"0001_00000_011_000", 	-- add a, r3
        42	=>	B"0110_00000_000_010", 	-- mov r2, a
        43	=>	B"0111_00000000000", 	-- clr c
        44	=>	B"0010_00000_101_000", 	-- subb a, r5
        45	=>	B"1110_000_11011111", 	-- jc loop
        46	=>	B"0101_00000010_010", 	-- mov r2, #2
        47	=>	B"0101_00000000_101", 	-- mov r5, #0
        48	=>	B"1001_00000_010_000", 	-- mov a, @r2
        49	=>	B"0110_00000_000_100", 	-- mov r4, a
        50	=>	B"1000_00000000_000", 	-- mov a, #0
        51	=>	B"0111_00000000000", 	-- clr c
        52	=>	B"0010_00000_100_000", 	-- subb a, r4
        53	=>	B"1110_000_00000111", 	-- jc mostrar
        54	=>	B"0001_00000_010_000", 	-- add a, r2
        55	=>	B"0001_00000_011_000", 	-- add a, r3
        56	=>	B"0110_00000_000_010", 	-- mov r2, a
        57	=>	B"0111_00000000000", 	-- clr c
        58	=>	B"0010_00000_001_000", 	-- subb a, r1
        59	=>	B"1110_000_11110100", 	-- jc ler_ram
        60	=>	B"1111_000_01000111", 	-- ajmp fim_leitura
        61	=>	B"1000_00000000_000", 	-- mov a, #0
        62	=>	B"0001_00000_100_000", 	-- add a, r4
        63	=>	B"0110_00000_000_101", 	-- mov r5, a
        64	=>	B"1000_00000000_000", 	-- mov a, #0
        65	=>	B"0001_00000_010_000", 	-- add a, r2
        66	=>	B"0001_00000_011_000", 	-- add a, r3
        67	=>	B"0110_00000_000_010", 	-- mov r2, a
        68	=>	B"0111_00000000000", 	-- clr c
        69	=>	B"0010_00000_001_000", 	-- subb a, r1
        70	=>	B"1110_000_11101001", 	-- jc ler_ram
        71	=>	B"0000_00000000000", 	-- nop

        others => (others=>'0')
    );

begin

    process(clk)
    begin
        if(rising_edge(clk)) then
            data <= conteudo_rom(to_integer(addr));
        end if;
    end process;
    
end architecture;