library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ula is
    port (
        clk : in std_logic;
        rst : in std_logic;
        sig
    );
end ula;

architecture rtl of a_ula is

begin

end architecture;